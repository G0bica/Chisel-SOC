module APBInterconnect(
  input         clock,
  input         reset,
  input  [31:0] io_in_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_in_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_in_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_in_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_in_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_in_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_in_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_in_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_0_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_0_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_0_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_0_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_0_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_0_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_0_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_0_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_1_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_1_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_1_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_1_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_1_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_1_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_1_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_1_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_2_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_2_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_2_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_2_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_2_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_2_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_2_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_2_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_3_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_3_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_3_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_3_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_3_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_3_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_3_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_3_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_4_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_4_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_4_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_4_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_4_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_4_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_4_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_4_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_5_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_5_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_5_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_5_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_5_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_5_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_5_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_5_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_6_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_6_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_6_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_6_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_6_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_6_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_6_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_6_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_7_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_7_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_7_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_7_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_7_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_7_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_7_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_7_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_8_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_8_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_8_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_8_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_8_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_8_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_8_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_8_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_9_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_9_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_9_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_9_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_9_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_9_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_9_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_9_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_10_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_10_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_10_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_10_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_10_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_10_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_10_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_10_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_11_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_11_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_11_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_11_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_11_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_11_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_11_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_11_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_12_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_12_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_12_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_12_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_12_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_12_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_12_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_12_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_13_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_13_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_13_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_13_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_13_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_13_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_13_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_13_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_14_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_14_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_14_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_14_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_14_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_14_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_14_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_14_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_15_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_15_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_15_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_15_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_15_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_15_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_15_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_15_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_16_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_16_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_16_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_16_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_16_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_16_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_16_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_16_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_17_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_17_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_17_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_17_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_17_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_17_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_17_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_17_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_18_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_18_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_18_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_18_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_18_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_18_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_18_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_18_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_19_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_19_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_19_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_19_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_19_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_19_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_19_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_19_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_20_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_20_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_20_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_20_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_20_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_20_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_20_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_20_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_21_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_21_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_21_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_21_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_21_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_21_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_21_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_21_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_22_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_22_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_22_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_22_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_22_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_22_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_22_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_22_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_23_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_23_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_23_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_23_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_23_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_23_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_23_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_23_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_24_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_24_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_24_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_24_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_24_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_24_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_24_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_24_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_25_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_25_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_25_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_25_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_25_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_25_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_25_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_25_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_26_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_26_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_26_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_26_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_26_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_26_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_26_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_26_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_27_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_27_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_27_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_27_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_27_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_27_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_27_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_27_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_28_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_28_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_28_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_28_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_28_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_28_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_28_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_28_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_29_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_29_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_29_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_29_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_29_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_29_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_29_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_29_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_30_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_30_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_30_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_30_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_30_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_30_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_30_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_30_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_31_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_31_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_31_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_31_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_31_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_31_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_31_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_31_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_32_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_32_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_32_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_32_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_32_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_32_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_32_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_32_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_33_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_33_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_33_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_33_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_33_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_33_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_33_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_33_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_34_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_34_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_34_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_34_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_34_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_34_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_34_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_34_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_35_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_35_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_35_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_35_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_35_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_35_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_35_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_35_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_36_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_36_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_36_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_36_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_36_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_36_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_36_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_36_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_37_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_37_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_37_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_37_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_37_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_37_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_37_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_37_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_38_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_38_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_38_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_38_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_38_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_38_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_38_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_38_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_39_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_39_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_39_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_39_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_39_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_39_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_39_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_39_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_40_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_40_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_40_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_40_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_40_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_40_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_40_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_40_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_41_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_41_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_41_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_41_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_41_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_41_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_41_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_41_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_42_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_42_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_42_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_42_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_42_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_42_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_42_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_42_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_43_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_43_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_43_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_43_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_43_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_43_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_43_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_43_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_44_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_44_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_44_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_44_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_44_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_44_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_44_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_44_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_45_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_45_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_45_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_45_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_45_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_45_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_45_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_45_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_46_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_46_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_46_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_46_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_46_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_46_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_46_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_46_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_47_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_47_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_47_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_47_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_47_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_47_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_47_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_47_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_48_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_48_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_48_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_48_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_48_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_48_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_48_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_48_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_49_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_49_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_49_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_49_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_49_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_49_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_49_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_49_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_50_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_50_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_50_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_50_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_50_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_50_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_50_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_50_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_51_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_51_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_51_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_51_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_51_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_51_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_51_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_51_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_52_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_52_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_52_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_52_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_52_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_52_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_52_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_52_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_53_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_53_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_53_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_53_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_53_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_53_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_53_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_53_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_54_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_54_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_54_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_54_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_54_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_54_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_54_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_54_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_55_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_55_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_55_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_55_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_55_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_55_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_55_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_55_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_56_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_56_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_56_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_56_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_56_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_56_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_56_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_56_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_57_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_57_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_57_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_57_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_57_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_57_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_57_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_57_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_58_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_58_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_58_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_58_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_58_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_58_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_58_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_58_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_59_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_59_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_59_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_59_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_59_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_59_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_59_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_59_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_60_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_60_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_60_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_60_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_60_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_60_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_60_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_60_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_61_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_61_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_61_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_61_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_61_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_61_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_61_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_61_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_62_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_62_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_62_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_62_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_62_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_62_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_62_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_62_pslverr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_63_psel, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_63_paddr, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_63_penable, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output        io_slaves_63_pwrite, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  output [31:0] io_slaves_63_pwdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input  [31:0] io_slaves_63_prdata, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_63_pready, // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
  input         io_slaves_63_pslverr // @[\\src\\main\\scala\\ApbInterconnect.scala 11:14]
);
  wire [5:0] peripheralIndex = io_in_paddr[12:7]; // @[\\src\\main\\scala\\ApbInterconnect.scala 44:36]
  wire  _GEN_1 = 6'h1 == peripheralIndex ? io_slaves_1_pready : io_slaves_0_pready; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_2 = 6'h2 == peripheralIndex ? io_slaves_2_pready : _GEN_1; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_3 = 6'h3 == peripheralIndex ? io_slaves_3_pready : _GEN_2; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_4 = 6'h4 == peripheralIndex ? io_slaves_4_pready : _GEN_3; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_5 = 6'h5 == peripheralIndex ? io_slaves_5_pready : _GEN_4; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_6 = 6'h6 == peripheralIndex ? io_slaves_6_pready : _GEN_5; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_7 = 6'h7 == peripheralIndex ? io_slaves_7_pready : _GEN_6; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_8 = 6'h8 == peripheralIndex ? io_slaves_8_pready : _GEN_7; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_9 = 6'h9 == peripheralIndex ? io_slaves_9_pready : _GEN_8; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_10 = 6'ha == peripheralIndex ? io_slaves_10_pready : _GEN_9; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_11 = 6'hb == peripheralIndex ? io_slaves_11_pready : _GEN_10; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_12 = 6'hc == peripheralIndex ? io_slaves_12_pready : _GEN_11; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_13 = 6'hd == peripheralIndex ? io_slaves_13_pready : _GEN_12; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_14 = 6'he == peripheralIndex ? io_slaves_14_pready : _GEN_13; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_15 = 6'hf == peripheralIndex ? io_slaves_15_pready : _GEN_14; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_16 = 6'h10 == peripheralIndex ? io_slaves_16_pready : _GEN_15; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_17 = 6'h11 == peripheralIndex ? io_slaves_17_pready : _GEN_16; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_18 = 6'h12 == peripheralIndex ? io_slaves_18_pready : _GEN_17; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_19 = 6'h13 == peripheralIndex ? io_slaves_19_pready : _GEN_18; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_20 = 6'h14 == peripheralIndex ? io_slaves_20_pready : _GEN_19; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_21 = 6'h15 == peripheralIndex ? io_slaves_21_pready : _GEN_20; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_22 = 6'h16 == peripheralIndex ? io_slaves_22_pready : _GEN_21; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_23 = 6'h17 == peripheralIndex ? io_slaves_23_pready : _GEN_22; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_24 = 6'h18 == peripheralIndex ? io_slaves_24_pready : _GEN_23; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_25 = 6'h19 == peripheralIndex ? io_slaves_25_pready : _GEN_24; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_26 = 6'h1a == peripheralIndex ? io_slaves_26_pready : _GEN_25; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_27 = 6'h1b == peripheralIndex ? io_slaves_27_pready : _GEN_26; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_28 = 6'h1c == peripheralIndex ? io_slaves_28_pready : _GEN_27; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_29 = 6'h1d == peripheralIndex ? io_slaves_29_pready : _GEN_28; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_30 = 6'h1e == peripheralIndex ? io_slaves_30_pready : _GEN_29; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_31 = 6'h1f == peripheralIndex ? io_slaves_31_pready : _GEN_30; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_32 = 6'h20 == peripheralIndex ? io_slaves_32_pready : _GEN_31; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_33 = 6'h21 == peripheralIndex ? io_slaves_33_pready : _GEN_32; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_34 = 6'h22 == peripheralIndex ? io_slaves_34_pready : _GEN_33; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_35 = 6'h23 == peripheralIndex ? io_slaves_35_pready : _GEN_34; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_36 = 6'h24 == peripheralIndex ? io_slaves_36_pready : _GEN_35; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_37 = 6'h25 == peripheralIndex ? io_slaves_37_pready : _GEN_36; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_38 = 6'h26 == peripheralIndex ? io_slaves_38_pready : _GEN_37; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_39 = 6'h27 == peripheralIndex ? io_slaves_39_pready : _GEN_38; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_40 = 6'h28 == peripheralIndex ? io_slaves_40_pready : _GEN_39; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_41 = 6'h29 == peripheralIndex ? io_slaves_41_pready : _GEN_40; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_42 = 6'h2a == peripheralIndex ? io_slaves_42_pready : _GEN_41; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_43 = 6'h2b == peripheralIndex ? io_slaves_43_pready : _GEN_42; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_44 = 6'h2c == peripheralIndex ? io_slaves_44_pready : _GEN_43; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_45 = 6'h2d == peripheralIndex ? io_slaves_45_pready : _GEN_44; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_46 = 6'h2e == peripheralIndex ? io_slaves_46_pready : _GEN_45; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_47 = 6'h2f == peripheralIndex ? io_slaves_47_pready : _GEN_46; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_48 = 6'h30 == peripheralIndex ? io_slaves_48_pready : _GEN_47; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_49 = 6'h31 == peripheralIndex ? io_slaves_49_pready : _GEN_48; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_50 = 6'h32 == peripheralIndex ? io_slaves_50_pready : _GEN_49; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_51 = 6'h33 == peripheralIndex ? io_slaves_51_pready : _GEN_50; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_52 = 6'h34 == peripheralIndex ? io_slaves_52_pready : _GEN_51; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_53 = 6'h35 == peripheralIndex ? io_slaves_53_pready : _GEN_52; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_54 = 6'h36 == peripheralIndex ? io_slaves_54_pready : _GEN_53; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_55 = 6'h37 == peripheralIndex ? io_slaves_55_pready : _GEN_54; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_56 = 6'h38 == peripheralIndex ? io_slaves_56_pready : _GEN_55; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_57 = 6'h39 == peripheralIndex ? io_slaves_57_pready : _GEN_56; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_58 = 6'h3a == peripheralIndex ? io_slaves_58_pready : _GEN_57; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_59 = 6'h3b == peripheralIndex ? io_slaves_59_pready : _GEN_58; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_60 = 6'h3c == peripheralIndex ? io_slaves_60_pready : _GEN_59; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_61 = 6'h3d == peripheralIndex ? io_slaves_61_pready : _GEN_60; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_62 = 6'h3e == peripheralIndex ? io_slaves_62_pready : _GEN_61; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  wire  _GEN_65 = 6'h1 == peripheralIndex ? io_slaves_1_pslverr : io_slaves_0_pslverr; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_66 = 6'h2 == peripheralIndex ? io_slaves_2_pslverr : _GEN_65; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_67 = 6'h3 == peripheralIndex ? io_slaves_3_pslverr : _GEN_66; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_68 = 6'h4 == peripheralIndex ? io_slaves_4_pslverr : _GEN_67; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_69 = 6'h5 == peripheralIndex ? io_slaves_5_pslverr : _GEN_68; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_70 = 6'h6 == peripheralIndex ? io_slaves_6_pslverr : _GEN_69; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_71 = 6'h7 == peripheralIndex ? io_slaves_7_pslverr : _GEN_70; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_72 = 6'h8 == peripheralIndex ? io_slaves_8_pslverr : _GEN_71; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_73 = 6'h9 == peripheralIndex ? io_slaves_9_pslverr : _GEN_72; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_74 = 6'ha == peripheralIndex ? io_slaves_10_pslverr : _GEN_73; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_75 = 6'hb == peripheralIndex ? io_slaves_11_pslverr : _GEN_74; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_76 = 6'hc == peripheralIndex ? io_slaves_12_pslverr : _GEN_75; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_77 = 6'hd == peripheralIndex ? io_slaves_13_pslverr : _GEN_76; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_78 = 6'he == peripheralIndex ? io_slaves_14_pslverr : _GEN_77; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_79 = 6'hf == peripheralIndex ? io_slaves_15_pslverr : _GEN_78; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_80 = 6'h10 == peripheralIndex ? io_slaves_16_pslverr : _GEN_79; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_81 = 6'h11 == peripheralIndex ? io_slaves_17_pslverr : _GEN_80; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_82 = 6'h12 == peripheralIndex ? io_slaves_18_pslverr : _GEN_81; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_83 = 6'h13 == peripheralIndex ? io_slaves_19_pslverr : _GEN_82; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_84 = 6'h14 == peripheralIndex ? io_slaves_20_pslverr : _GEN_83; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_85 = 6'h15 == peripheralIndex ? io_slaves_21_pslverr : _GEN_84; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_86 = 6'h16 == peripheralIndex ? io_slaves_22_pslverr : _GEN_85; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_87 = 6'h17 == peripheralIndex ? io_slaves_23_pslverr : _GEN_86; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_88 = 6'h18 == peripheralIndex ? io_slaves_24_pslverr : _GEN_87; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_89 = 6'h19 == peripheralIndex ? io_slaves_25_pslverr : _GEN_88; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_90 = 6'h1a == peripheralIndex ? io_slaves_26_pslverr : _GEN_89; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_91 = 6'h1b == peripheralIndex ? io_slaves_27_pslverr : _GEN_90; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_92 = 6'h1c == peripheralIndex ? io_slaves_28_pslverr : _GEN_91; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_93 = 6'h1d == peripheralIndex ? io_slaves_29_pslverr : _GEN_92; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_94 = 6'h1e == peripheralIndex ? io_slaves_30_pslverr : _GEN_93; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_95 = 6'h1f == peripheralIndex ? io_slaves_31_pslverr : _GEN_94; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_96 = 6'h20 == peripheralIndex ? io_slaves_32_pslverr : _GEN_95; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_97 = 6'h21 == peripheralIndex ? io_slaves_33_pslverr : _GEN_96; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_98 = 6'h22 == peripheralIndex ? io_slaves_34_pslverr : _GEN_97; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_99 = 6'h23 == peripheralIndex ? io_slaves_35_pslverr : _GEN_98; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_100 = 6'h24 == peripheralIndex ? io_slaves_36_pslverr : _GEN_99; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_101 = 6'h25 == peripheralIndex ? io_slaves_37_pslverr : _GEN_100; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_102 = 6'h26 == peripheralIndex ? io_slaves_38_pslverr : _GEN_101; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_103 = 6'h27 == peripheralIndex ? io_slaves_39_pslverr : _GEN_102; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_104 = 6'h28 == peripheralIndex ? io_slaves_40_pslverr : _GEN_103; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_105 = 6'h29 == peripheralIndex ? io_slaves_41_pslverr : _GEN_104; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_106 = 6'h2a == peripheralIndex ? io_slaves_42_pslverr : _GEN_105; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_107 = 6'h2b == peripheralIndex ? io_slaves_43_pslverr : _GEN_106; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_108 = 6'h2c == peripheralIndex ? io_slaves_44_pslverr : _GEN_107; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_109 = 6'h2d == peripheralIndex ? io_slaves_45_pslverr : _GEN_108; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_110 = 6'h2e == peripheralIndex ? io_slaves_46_pslverr : _GEN_109; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_111 = 6'h2f == peripheralIndex ? io_slaves_47_pslverr : _GEN_110; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_112 = 6'h30 == peripheralIndex ? io_slaves_48_pslverr : _GEN_111; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_113 = 6'h31 == peripheralIndex ? io_slaves_49_pslverr : _GEN_112; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_114 = 6'h32 == peripheralIndex ? io_slaves_50_pslverr : _GEN_113; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_115 = 6'h33 == peripheralIndex ? io_slaves_51_pslverr : _GEN_114; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_116 = 6'h34 == peripheralIndex ? io_slaves_52_pslverr : _GEN_115; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_117 = 6'h35 == peripheralIndex ? io_slaves_53_pslverr : _GEN_116; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_118 = 6'h36 == peripheralIndex ? io_slaves_54_pslverr : _GEN_117; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_119 = 6'h37 == peripheralIndex ? io_slaves_55_pslverr : _GEN_118; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_120 = 6'h38 == peripheralIndex ? io_slaves_56_pslverr : _GEN_119; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_121 = 6'h39 == peripheralIndex ? io_slaves_57_pslverr : _GEN_120; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_122 = 6'h3a == peripheralIndex ? io_slaves_58_pslverr : _GEN_121; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_123 = 6'h3b == peripheralIndex ? io_slaves_59_pslverr : _GEN_122; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_124 = 6'h3c == peripheralIndex ? io_slaves_60_pslverr : _GEN_123; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_125 = 6'h3d == peripheralIndex ? io_slaves_61_pslverr : _GEN_124; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire  _GEN_126 = 6'h3e == peripheralIndex ? io_slaves_62_pslverr : _GEN_125; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  wire [31:0] _GEN_129 = 6'h1 == peripheralIndex ? io_slaves_1_prdata : io_slaves_0_prdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_130 = 6'h2 == peripheralIndex ? io_slaves_2_prdata : _GEN_129; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_131 = 6'h3 == peripheralIndex ? io_slaves_3_prdata : _GEN_130; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_132 = 6'h4 == peripheralIndex ? io_slaves_4_prdata : _GEN_131; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_133 = 6'h5 == peripheralIndex ? io_slaves_5_prdata : _GEN_132; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_134 = 6'h6 == peripheralIndex ? io_slaves_6_prdata : _GEN_133; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_135 = 6'h7 == peripheralIndex ? io_slaves_7_prdata : _GEN_134; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_136 = 6'h8 == peripheralIndex ? io_slaves_8_prdata : _GEN_135; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_137 = 6'h9 == peripheralIndex ? io_slaves_9_prdata : _GEN_136; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_138 = 6'ha == peripheralIndex ? io_slaves_10_prdata : _GEN_137; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_139 = 6'hb == peripheralIndex ? io_slaves_11_prdata : _GEN_138; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_140 = 6'hc == peripheralIndex ? io_slaves_12_prdata : _GEN_139; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_141 = 6'hd == peripheralIndex ? io_slaves_13_prdata : _GEN_140; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_142 = 6'he == peripheralIndex ? io_slaves_14_prdata : _GEN_141; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_143 = 6'hf == peripheralIndex ? io_slaves_15_prdata : _GEN_142; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_144 = 6'h10 == peripheralIndex ? io_slaves_16_prdata : _GEN_143; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_145 = 6'h11 == peripheralIndex ? io_slaves_17_prdata : _GEN_144; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_146 = 6'h12 == peripheralIndex ? io_slaves_18_prdata : _GEN_145; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_147 = 6'h13 == peripheralIndex ? io_slaves_19_prdata : _GEN_146; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_148 = 6'h14 == peripheralIndex ? io_slaves_20_prdata : _GEN_147; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_149 = 6'h15 == peripheralIndex ? io_slaves_21_prdata : _GEN_148; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_150 = 6'h16 == peripheralIndex ? io_slaves_22_prdata : _GEN_149; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_151 = 6'h17 == peripheralIndex ? io_slaves_23_prdata : _GEN_150; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_152 = 6'h18 == peripheralIndex ? io_slaves_24_prdata : _GEN_151; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_153 = 6'h19 == peripheralIndex ? io_slaves_25_prdata : _GEN_152; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_154 = 6'h1a == peripheralIndex ? io_slaves_26_prdata : _GEN_153; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_155 = 6'h1b == peripheralIndex ? io_slaves_27_prdata : _GEN_154; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_156 = 6'h1c == peripheralIndex ? io_slaves_28_prdata : _GEN_155; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_157 = 6'h1d == peripheralIndex ? io_slaves_29_prdata : _GEN_156; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_158 = 6'h1e == peripheralIndex ? io_slaves_30_prdata : _GEN_157; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_159 = 6'h1f == peripheralIndex ? io_slaves_31_prdata : _GEN_158; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_160 = 6'h20 == peripheralIndex ? io_slaves_32_prdata : _GEN_159; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_161 = 6'h21 == peripheralIndex ? io_slaves_33_prdata : _GEN_160; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_162 = 6'h22 == peripheralIndex ? io_slaves_34_prdata : _GEN_161; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_163 = 6'h23 == peripheralIndex ? io_slaves_35_prdata : _GEN_162; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_164 = 6'h24 == peripheralIndex ? io_slaves_36_prdata : _GEN_163; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_165 = 6'h25 == peripheralIndex ? io_slaves_37_prdata : _GEN_164; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_166 = 6'h26 == peripheralIndex ? io_slaves_38_prdata : _GEN_165; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_167 = 6'h27 == peripheralIndex ? io_slaves_39_prdata : _GEN_166; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_168 = 6'h28 == peripheralIndex ? io_slaves_40_prdata : _GEN_167; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_169 = 6'h29 == peripheralIndex ? io_slaves_41_prdata : _GEN_168; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_170 = 6'h2a == peripheralIndex ? io_slaves_42_prdata : _GEN_169; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_171 = 6'h2b == peripheralIndex ? io_slaves_43_prdata : _GEN_170; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_172 = 6'h2c == peripheralIndex ? io_slaves_44_prdata : _GEN_171; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_173 = 6'h2d == peripheralIndex ? io_slaves_45_prdata : _GEN_172; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_174 = 6'h2e == peripheralIndex ? io_slaves_46_prdata : _GEN_173; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_175 = 6'h2f == peripheralIndex ? io_slaves_47_prdata : _GEN_174; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_176 = 6'h30 == peripheralIndex ? io_slaves_48_prdata : _GEN_175; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_177 = 6'h31 == peripheralIndex ? io_slaves_49_prdata : _GEN_176; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_178 = 6'h32 == peripheralIndex ? io_slaves_50_prdata : _GEN_177; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_179 = 6'h33 == peripheralIndex ? io_slaves_51_prdata : _GEN_178; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_180 = 6'h34 == peripheralIndex ? io_slaves_52_prdata : _GEN_179; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_181 = 6'h35 == peripheralIndex ? io_slaves_53_prdata : _GEN_180; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_182 = 6'h36 == peripheralIndex ? io_slaves_54_prdata : _GEN_181; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_183 = 6'h37 == peripheralIndex ? io_slaves_55_prdata : _GEN_182; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_184 = 6'h38 == peripheralIndex ? io_slaves_56_prdata : _GEN_183; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_185 = 6'h39 == peripheralIndex ? io_slaves_57_prdata : _GEN_184; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_186 = 6'h3a == peripheralIndex ? io_slaves_58_prdata : _GEN_185; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_187 = 6'h3b == peripheralIndex ? io_slaves_59_prdata : _GEN_186; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_188 = 6'h3c == peripheralIndex ? io_slaves_60_prdata : _GEN_187; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_189 = 6'h3d == peripheralIndex ? io_slaves_61_prdata : _GEN_188; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_190 = 6'h3e == peripheralIndex ? io_slaves_62_prdata : _GEN_189; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  wire [31:0] _GEN_191 = 6'h3f == peripheralIndex ? io_slaves_63_prdata : _GEN_190; // @[\\src\\main\\scala\\ApbInterconnect.scala 66:{18,18}]
  assign io_in_prdata = ~io_in_pwrite & io_in_psel ? _GEN_191 : 32'h0; // @[\\src\\main\\scala\\ApbInterconnect.scala 64:16 65:37 66:18]
  assign io_in_pready = 6'h3f == peripheralIndex ? io_slaves_63_pready : _GEN_62; // @[\\src\\main\\scala\\ApbInterconnect.scala 60:{17,17}]
  assign io_in_pslverr = 6'h3f == peripheralIndex ? io_slaves_63_pslverr : _GEN_126; // @[\\src\\main\\scala\\ApbInterconnect.scala 61:{17,17}]
  assign io_slaves_0_psel = io_in_psel & peripheralIndex == 6'h0; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_0_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_0_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_0_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_0_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_1_psel = io_in_psel & peripheralIndex == 6'h1; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_1_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_1_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_1_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_1_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_2_psel = io_in_psel & peripheralIndex == 6'h2; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_2_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_2_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_2_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_2_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_3_psel = io_in_psel & peripheralIndex == 6'h3; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_3_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_3_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_3_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_3_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_4_psel = io_in_psel & peripheralIndex == 6'h4; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_4_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_4_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_4_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_4_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_5_psel = io_in_psel & peripheralIndex == 6'h5; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_5_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_5_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_5_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_5_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_6_psel = io_in_psel & peripheralIndex == 6'h6; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_6_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_6_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_6_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_6_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_7_psel = io_in_psel & peripheralIndex == 6'h7; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_7_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_7_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_7_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_7_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_8_psel = io_in_psel & peripheralIndex == 6'h8; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_8_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_8_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_8_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_8_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_9_psel = io_in_psel & peripheralIndex == 6'h9; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_9_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_9_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_9_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_9_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_10_psel = io_in_psel & peripheralIndex == 6'ha; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_10_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_10_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_10_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_10_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_11_psel = io_in_psel & peripheralIndex == 6'hb; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_11_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_11_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_11_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_11_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_12_psel = io_in_psel & peripheralIndex == 6'hc; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_12_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_12_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_12_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_12_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_13_psel = io_in_psel & peripheralIndex == 6'hd; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_13_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_13_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_13_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_13_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_14_psel = io_in_psel & peripheralIndex == 6'he; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_14_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_14_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_14_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_14_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_15_psel = io_in_psel & peripheralIndex == 6'hf; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_15_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_15_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_15_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_15_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_16_psel = io_in_psel & peripheralIndex == 6'h10; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_16_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_16_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_16_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_16_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_17_psel = io_in_psel & peripheralIndex == 6'h11; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_17_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_17_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_17_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_17_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_18_psel = io_in_psel & peripheralIndex == 6'h12; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_18_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_18_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_18_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_18_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_19_psel = io_in_psel & peripheralIndex == 6'h13; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_19_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_19_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_19_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_19_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_20_psel = io_in_psel & peripheralIndex == 6'h14; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_20_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_20_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_20_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_20_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_21_psel = io_in_psel & peripheralIndex == 6'h15; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_21_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_21_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_21_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_21_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_22_psel = io_in_psel & peripheralIndex == 6'h16; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_22_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_22_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_22_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_22_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_23_psel = io_in_psel & peripheralIndex == 6'h17; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_23_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_23_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_23_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_23_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_24_psel = io_in_psel & peripheralIndex == 6'h18; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_24_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_24_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_24_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_24_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_25_psel = io_in_psel & peripheralIndex == 6'h19; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_25_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_25_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_25_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_25_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_26_psel = io_in_psel & peripheralIndex == 6'h1a; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_26_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_26_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_26_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_26_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_27_psel = io_in_psel & peripheralIndex == 6'h1b; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_27_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_27_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_27_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_27_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_28_psel = io_in_psel & peripheralIndex == 6'h1c; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_28_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_28_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_28_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_28_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_29_psel = io_in_psel & peripheralIndex == 6'h1d; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_29_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_29_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_29_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_29_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_30_psel = io_in_psel & peripheralIndex == 6'h1e; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_30_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_30_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_30_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_30_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_31_psel = io_in_psel & peripheralIndex == 6'h1f; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_31_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_31_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_31_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_31_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_32_psel = io_in_psel & peripheralIndex == 6'h20; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_32_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_32_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_32_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_32_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_33_psel = io_in_psel & peripheralIndex == 6'h21; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_33_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_33_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_33_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_33_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_34_psel = io_in_psel & peripheralIndex == 6'h22; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_34_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_34_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_34_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_34_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_35_psel = io_in_psel & peripheralIndex == 6'h23; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_35_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_35_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_35_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_35_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_36_psel = io_in_psel & peripheralIndex == 6'h24; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_36_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_36_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_36_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_36_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_37_psel = io_in_psel & peripheralIndex == 6'h25; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_37_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_37_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_37_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_37_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_38_psel = io_in_psel & peripheralIndex == 6'h26; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_38_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_38_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_38_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_38_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_39_psel = io_in_psel & peripheralIndex == 6'h27; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_39_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_39_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_39_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_39_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_40_psel = io_in_psel & peripheralIndex == 6'h28; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_40_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_40_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_40_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_40_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_41_psel = io_in_psel & peripheralIndex == 6'h29; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_41_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_41_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_41_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_41_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_42_psel = io_in_psel & peripheralIndex == 6'h2a; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_42_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_42_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_42_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_42_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_43_psel = io_in_psel & peripheralIndex == 6'h2b; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_43_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_43_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_43_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_43_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_44_psel = io_in_psel & peripheralIndex == 6'h2c; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_44_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_44_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_44_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_44_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_45_psel = io_in_psel & peripheralIndex == 6'h2d; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_45_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_45_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_45_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_45_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_46_psel = io_in_psel & peripheralIndex == 6'h2e; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_46_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_46_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_46_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_46_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_47_psel = io_in_psel & peripheralIndex == 6'h2f; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_47_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_47_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_47_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_47_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_48_psel = io_in_psel & peripheralIndex == 6'h30; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_48_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_48_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_48_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_48_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_49_psel = io_in_psel & peripheralIndex == 6'h31; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_49_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_49_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_49_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_49_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_50_psel = io_in_psel & peripheralIndex == 6'h32; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_50_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_50_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_50_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_50_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_51_psel = io_in_psel & peripheralIndex == 6'h33; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_51_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_51_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_51_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_51_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_52_psel = io_in_psel & peripheralIndex == 6'h34; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_52_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_52_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_52_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_52_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_53_psel = io_in_psel & peripheralIndex == 6'h35; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_53_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_53_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_53_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_53_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_54_psel = io_in_psel & peripheralIndex == 6'h36; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_54_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_54_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_54_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_54_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_55_psel = io_in_psel & peripheralIndex == 6'h37; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_55_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_55_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_55_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_55_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_56_psel = io_in_psel & peripheralIndex == 6'h38; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_56_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_56_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_56_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_56_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_57_psel = io_in_psel & peripheralIndex == 6'h39; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_57_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_57_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_57_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_57_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_58_psel = io_in_psel & peripheralIndex == 6'h3a; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_58_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_58_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_58_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_58_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_59_psel = io_in_psel & peripheralIndex == 6'h3b; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_59_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_59_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_59_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_59_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_60_psel = io_in_psel & peripheralIndex == 6'h3c; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_60_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_60_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_60_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_60_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_61_psel = io_in_psel & peripheralIndex == 6'h3d; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_61_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_61_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_61_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_61_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_62_psel = io_in_psel & peripheralIndex == 6'h3e; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_62_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_62_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_62_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_62_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
  assign io_slaves_63_psel = io_in_psel & peripheralIndex == 6'h3f; // @[\\src\\main\\scala\\ApbInterconnect.scala 55:37]
  assign io_slaves_63_paddr = io_in_paddr; // @[\\src\\main\\scala\\ApbInterconnect.scala 49:26]
  assign io_slaves_63_penable = io_in_penable; // @[\\src\\main\\scala\\ApbInterconnect.scala 50:26]
  assign io_slaves_63_pwrite = io_in_pwrite; // @[\\src\\main\\scala\\ApbInterconnect.scala 51:26]
  assign io_slaves_63_pwdata = io_in_pwdata; // @[\\src\\main\\scala\\ApbInterconnect.scala 52:26]
endmodule
